`include "../../lib/EECS151.v"

module structural_adder #(
    parameter N = 3
) (
    input [N-1:0] a,
    input [N-1:0] b,
    output [N:0] sum
);
    // TODO: Your code (from lab 2). You need to parameterize it

endmodule

`timescale 1ns/1ns

// UART_Transmitter is essentially a reverse of UART_Receiver
module uart_transmitter_tb();
    localparam CLOCK_FREQUENCY  = 125_000_000;
    localparam CLOCK_PERIOD     = 1_000_000_000 / CLOCK_FREQUENCY;
    localparam BAUD_RATE        = 115_200;
    localparam BAUD_PERIOD      = 1_000_000_000 / BAUD_RATE; // 8680.55 ns

    localparam CHAR0 = 8'h61; // ~ 'a'
    localparam NUM_CHARS = 10;

    reg clk, rst;
    initial clk = 0;
    always #(CLOCK_PERIOD / 2) clk = ~clk;
    
    wire [7:0] data_in;
    reg data_in_valid;
    wire data_in_ready;
    wire serial_out;

    uart_transmitter #(
        .CLOCK_FREQ(CLOCK_FREQUENCY),
        .BAUD_RATE(BAUD_RATE)
    ) dut (
        .clk(clk),
        .rst(rst),

        .data_in(data_in),             // input
        .data_in_valid(data_in_valid), // input
        .data_in_ready(data_in_ready), // output
        .serial_out(serial_out)        // output
    );

    reg data_in_fired;
    integer i, c;

    // this holds characters sent by the UART_transmitter to the host via serial line
    // including the start and stop bits
    reg [10-1:0] chars_to_host [NUM_CHARS-1:0];
    // this holds characters to be enqueued to data_in via R/V
    reg [7:0] chars_from_data_in [NUM_CHARS-1:0];

    // initialize test vectors
    initial begin
        #0
        for (c = 0; c < NUM_CHARS; c = c + 1) begin
           chars_from_data_in[c] = CHAR0 + c;
        end
    end

    reg [31:0] cnt;

    assign data_in = chars_from_data_in[cnt];

    always @(posedge clk) begin
        // data considered "enqueued" ("fired") when both valid and ready are
        // HIGH
        if (data_in_valid & data_in_ready) begin
            data_in_fired <= 1'b1;
            cnt <= cnt + 1;
            $display("[time %t] [data_in] Sent char: 8'h%h", $time, data_in);
        end

        // Set data_in_valid to LOW after we have sent all characters
        if (cnt == NUM_CHARS)
            data_in_valid <= 1'b0;

        // data_in_ready should be LOW in the next rising edge
        // after "fired"
        if (data_in_fired) begin
            if (data_in_ready == 1'b1) begin
                $display("[time %t] Failed: data_in_ready should go LOW after firing data_in\n", $time);
                $finish();
            end
            data_in_fired <= 1'b0;
        end
    end

    integer num_mismatches = 0;

    initial begin
        #0;
        rst = 1;
        data_in_valid = 0;
        cnt = 0;

        // Hold reset for a while
        repeat (10) @(posedge clk);

        rst = 0;

        if (data_in_ready == 1'b0) begin
            $display("[time %t] Failed: data_in_ready should not be LOW initially", $time);
            $finish();
        end

        // Delay for some time
        repeat (100) @(posedge clk);

        // The testbench has valid data to send to UART_Transmitter
        data_in_valid = 1;

        for (c = 0; c < NUM_CHARS; c = c + 1) begin
            // Wait until serial_out is LOW (start of transaction)
            while (serial_out == 1) begin
                @(posedge clk);
            end

            for (i = 0; i < 10; i = i + 1) begin
                chars_to_host[c][i] = serial_out;
                #(BAUD_PERIOD);
            end
            $display("[time %t] [serial_out] Got char: start_bit=%b, payload=8'h%h, stop_bit=%b", $time,
                chars_to_host[c][0], chars_to_host[c][8:1], chars_to_host[c][9]);
        end

        // Delay for some time
        repeat (10) @(posedge clk);

        // Check results
        for (c = 0; c < NUM_CHARS; c = c + 1) begin
            if (chars_from_data_in[c] !== chars_to_host[c][8:1]) begin
                $display("Mismatches at char %d: char_to_host=%h, char_from_data_in=%h",
                         c, chars_to_host[c], chars_from_data_in[c]);
                num_mismatches = num_mismatches + 1;
            end
            if (chars_to_host[c][0] != 0)
                $display("[char #%d] Failed: Start bit is not 0!", c);
            if (chars_to_host[c][9] != 1)
                $display("[char #%d] Failed: End bit is not 1!", c);
        end

        if (serial_out != 1) begin
            $display("Failed: serial_out should stay HIGH if there is no data_in to enqueue!");
            $finish();
        end

        $display("Test passed!");
        #100;
        $finish();
    end

    initial begin
        #(BAUD_PERIOD * 10 * (NUM_CHARS + 1));
        $display("TIMEOUT");
        $finish();
    end
endmodule

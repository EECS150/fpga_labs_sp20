`include "../../lib/EECS151.v"

module counter #(
    parameter N = 4,
    parameter RATE_HZ = 1
) (
    input clk,
    input rst_counter,
    input [N-1:0] rst_counter_val,
    output [N-1:0] counter_output
);

    //TODO : Your code

endmodule
